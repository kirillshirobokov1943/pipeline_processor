`include "defines.svh"
module instr_mem #(parameter width = 32, depth = 256)
(
	input logic                        arstn,
	input logic  [$clog2(depth)-1 : 0] A,
	output logic [width-1:0]           instr
);	
logic [width-1:0] data [depth-1:0];

//прошивка памяти инструкций при сбросе
always_ff @(negedge arstn) begin
//основной код для проверки - в под конец программы a0=2

data[0] <= 32'h00200613;
data[1] <= 32'h00300693;
data[2] <= 32'h00e00913;
data[3] <= 32'h00a00993;
data[4] <= 32'h00000393;
data[5] <= 32'h00000313;
data[6] <= 32'h00000413;
data[7] <= 32'h00c383b3;
data[8] <= 32'h00140413;
data[9] <= 32'hff241ce3;
data[10] <= 32'h00000413;
data[11] <= 32'h00d30333;
data[12] <= 32'h00140413;
data[13] <= 32'hff341ce3;
data[14] <= 32'h00100413;
data[15] <= 32'h40730533;
data[16] <= 32'hfc1ff7ef;
for (int i= 17; i<depth; i++)
   data[i] <= 32'd0;

    //код на проверку условных переходов назад
	 /*
   data[0] <= 32'h00000537;
	data[1] <= 32'h01e00613;
	
	data[2] <= 32'h00000593;
	
	data[3] <= 32'h01e58593;
	data[4] <= 32'h00a50513;
	data[5] <= 32'hfec58ce3;
	data[6] <= 32'h00700513;
	*/
	
	//код на проверку словных переходов вперед (с beq)
	/*
	data[0] <=32'h00000513 ;
	data[1] <=32'h00050863 ;
	data[2] <=32'h00700513 ;
	data[3] <=32'h00700513 ;
	data[4] <=32'h00700513 ;
	data[5] <=32'h00500513 ;
	data[6] <=32'h00800513 ;
	data[7] <=32'h00900513 ;
	data[8] <=32'h00400513 ;
	*/
	
	//код на проверку словных переходов вперед (с bne)
	/*
	data[0] <=32'h00300513 ;
	data[1] <=32'h00051863 ;
	data[2] <=32'h00700513 ;
	data[3] <=32'h00700513 ;
	data[4] <=32'h00600513 ;
	data[5] <=32'h00500513 ;
	data[6] <=32'h00800513 ;
	data[7] <=32'h00900513 ;
	*/
	
	
	//код на проверку безусловных переходов
	/*
	data[0] <=32'h00000513 ;
	data[1] <=32'h00c0056f ;
	data[2] <=32'h00100513 ;
	data[3] <=32'h00200513 ;
	data[4] <=32'h00300513 ;
	data[5] <=32'h00500513 ;
	*/
	
	
//случайная прорамма 1:
/*
data[0] <=32'h00001537;
data[1] <=32'h00550513;
data[2] <=32'h01400293;
data[3] <=32'h00550533;
data[4] <=32'h00f00313;
data[5] <=32'h00656533;
data[6] <=32'h00655533;
data[7] <=32'h40550533;
data[8] <=32'h00a00393;
data[9] <=32'h00753533;
data[10] <=32'h00500e13;
data[11] <=32'h00150513;
data[12] <=32'h00500e13;
data[13] <=32'h00750463;
data[14] <=32'hffc51ae3;
data[15] <=32'h048000ef;
data[16] <=32'h00150513;
data[17] <=32'h01d50533;
data[18] <=32'h03200e93;
data[19] <=32'h00a00513;
data[20] <=32'h41d50533;
data[21] <=32'h01d56533;
data[22] <=32'h01d55533;
data[23] <=32'h01d53533;
data[24] <=32'h00250513;
data[25] <=32'h00a50533;
data[26] <=32'h40a50533;
data[27] <=32'hf95ff96f;
data[28] <=32'h00a00f13;
data[29] <=32'h00350513;
data[30] <=32'h401f0f33;
data[31] <=32'hfe0f1ce3;
data[32] <=32'h00a00893;
data[33] <=32'h06450513;
data[34] <=32'h00556533;
data[35] <=32'h00655533;
data[36] <=32'h40750533;
data[37] <=32'h01c53533;
data[38] <=32'hfb1ff56f;
*/

  //слцчайная программа  2
/*
data[0] <= 32'h00000537;
data[1] <=32'h00050513;
data[2] <=32'h01900f93;
data[3] <=32'h00100293;
data[4] <=32'h00a00313;
data[5] <=32'h000283b3;
data[6] <=32'h00000e33;
data[7] <=32'h00028eb3;
data[8] <=32'h00750533;
data[9] <=32'hfffe8e93;
data[10] <=32'hfe0e9ce3;
data[11] <=32'h01c50533;
data[12] <=32'h01f50c63;
data[13] <=32'h00128293;
data[14] <=32'h00533533;
data[15] <=32'hfc050ce3;
data[16] <=32'h00656533;
data[17] <=32'h00555533;
data[18] <=32'h00656533;
data[19] <=32'h00550513;
data[20] <=32'h0180056f;
data[21] <=32'h00150513;
data[22] <=32'h00050463;
data[23] <=32'hfe051ce3;
data[24] <=32'h00a00893;
data[25] <=32'h00000073;
data[26] <=32'h06400513;
data[27] <=32'h00556533;
data[28] <=32'h00655533;
data[29] <=32'h40750533;
data[30] <=32'h01c53533;
data[31] <=32'hf85ff06f;
*/

     //тестовая программа 3
/*
data[0] <=32'hffc18537;
data[1] <=32'h00050513;
data[2] <=32'h00100293;
data[3] <=32'h00a00313;
data[4] <=32'h00100393;
data[5] <=32'h00039463;
data[6] <=32'h00550533;
data[7] <=32'h00130513;
data[8] <=32'h00533533;
data[9] <=32'h000e0463;
data[10] <=32'h00656533;
data[11] <=32'h00555533;
data[12] <=32'h40650533;
data[13] <=32'h00550513;
data[14] <=32'h0140006f;
data[15] <=32'h00150513;
data[16] <=32'h00050463;
data[17] <=32'hfe051ce3;
data[18] <=32'h00a00893;
data[19] <=32'h06450513;
data[20] <=32'h00556533;
data[21] <=32'h00655533;
data[22] <=32'h40750533;
data[23] <=32'h00a00e13;
data[24] <=32'h01c53533;
data[25] <=32'hfa1ff06f;
*/

    //тестовая программа 4
/*
data[0] <=32'h00000537;
data[1] <=32'h00750513;
data[2] <=32'h00300293;
data[3] <=32'h00f00313;
data[4] <=32'h00100393;
data[5] <=32'h00650533;
data[6] <=32'h40750533;
data[7] <=32'h00556533;
data[8] <=32'h00755533;
data[9] <=32'hfff28293;
data[10] <=32'hfe0296e3;
data[11] <=32'h03200e13;
data[12] <=32'h01c53eb3;
data[13] <=32'h000e8863;
data[14] <=32'h06450513;
data[15] <=32'h034000ef;
data[16] <=32'h0100006f;
data[17] <=32'h41c50533;
data[18] <=32'h01c56533;
data[19] <=32'h024000ef;
data[20] <=32'h00150513;
data[21] <=32'h00500f13;
data[22] <=32'h01e50533;
data[23] <=32'h40750533;
data[24] <=32'h00755533;
data[25] <=32'hffff0f13;
data[26] <=32'hfe0f18e3;
data[27] <=32'h00a00893;
data[28] <=32'h02a50513;
data[29] <=32'h00653533;
data[30] <=32'h00750533;
data[31] <=32'hf85ff06f;
*/



end	
	
logic [$clog2(depth)-1 : 0] addr;
assign addr = A>>2;
assign instr = data[addr];
endmodule